library work;
package Common is
  constant IPWM_DATA_WIDTH : integer := 8;

end Common;

package body Common is
  -- subprogram bodies here
end Common;