----------------------------------------------------------------------------
--	btn_debounce_toggle.vhd -- Button Debouncer
----------------------------------------------------------------------------
-- Author:  Sam Bobrowicz
--          Copyright 2011 Digilent, Inc.
-- Modified: Added toggle output
----------------------------------------------------------------------------
--
----------------------------------------------------------------------------
-- This component is used to debounce signals generated by external push
-- buttons. It is designed to independently debounce a Push button signal.
-- Debouncing is done by only registering a change in a button state if 
-- it remains constant for 2^16 clock cycles. 
--         				
-- Port Descriptions:
--
--   BTN_I 		- The input button signals
--   CLK  		- Behavior is optimized for a 100 MHz clock
--   BTN_O 		- The debounced button signals
--   TOGGLE_O 	- Debounced toggle output										
----------------------------------------------------------------------------
--
----------------------------------------------------------------------------
-- Revision History:
--  08/08/2011(SamB): Created using Xilinx Tools 13.2
--  10/06/2013  (CU): Converted to one button and added toggle output
----------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_unsigned.all;

entity btn_debounce_toggle is
GENERIC (
	CONSTANT CNTR_MAX : std_logic_vector(15 downto 0) := X"FFFF");
    Port ( BTN_I 	: in  STD_LOGIC;
           CLK 		: in  STD_LOGIC;
           BTN_O 	: out  STD_LOGIC;
			  pulse_O :out std_logic;
           TOGGLE_O : out  STD_LOGIC);
end btn_debounce_toggle;

architecture Behavioral of btn_debounce_toggle is

--constant CNTR_MAX : std_logic_vector(15 downto 0) := X"1";
signal btn_cntr   : std_logic_vector(15 downto 0) := (others => '0');
signal btn_reg    : std_logic   				  := '0';
signal btn_toggle : std_logic                     := '0';
signal btn_sync   : std_logic_vector(1 downto 0)  := (others => '1');
signal btn_pulse  : std_logic                     := '0';
signal btn_pulse_f: std_logic							  := '0';


begin

	btn_debounce_process : process (CLK)
	begin
		if (rising_edge(CLK)) then
			if (btn_cntr = CNTR_MAX) then
				btn_reg <= not(btn_reg);
			end if;
		end if;
	end process;
	
	btn_counter_process : process (CLK)
	begin
		if (rising_edge(CLK)) then
			if ((btn_reg = '1') xor (BTN_I = '1')) then
				if (btn_cntr = CNTR_MAX) then
					btn_cntr <= (others => '0');
				else
					btn_cntr <= btn_cntr + 1;
				end if;
			else
				btn_cntr <= (others => '0');
			end if;
		end if;
	end process;
	
	btn_toggle_process : process(CLK)
	begin
		if (rising_edge(CLK)) then
			btn_sync(0) <= btn_reg;
			btn_sync(1) <= btn_sync(0);
			btn_pulse   <= not btn_sync(1) and btn_sync(0);	--rising  edge
			btn_pulse_f <= btn_sync(1) and not btn_sync(0);	--falling edge
				if 	btn_pulse = '1' then
					btn_toggle <= not btn_toggle;
				end if;
		end if;
	end process;
					  
	BTN_O <= btn_reg;
	TOGGLE_O <= btn_toggle;
	pulse_O <= btn_pulse_f;

end Behavioral;